
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_test_state_buffer.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_test_state_buffer.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_test_state_buffer.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_34_1_fu_7484.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_34_1_fu_7484.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_34_1_fu_7484.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_39_2_fu_7490.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_39_2_fu_7490.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_39_2_fu_7490.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;

    seq_loop_intf#(276) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state5;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state265;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state263;
    assign seq_loop_intf_1.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.quit_loop_state1 = AESL_inst_test_state_buffer.ap_ST_fsm_state264;
    assign seq_loop_intf_1.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state262;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state264;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(276) seq_loop_monitor_1;
    seq_loop_intf#(276) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state5;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state9;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state8;
    assign seq_loop_intf_2.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_2.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state6;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state8;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(276) seq_loop_monitor_2;
    seq_loop_intf#(276) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state9;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state13;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state12;
    assign seq_loop_intf_3.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_3.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state10;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state12;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(276) seq_loop_monitor_3;
    seq_loop_intf#(276) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state13;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state17;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state16;
    assign seq_loop_intf_4.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_4.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state14;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state16;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(276) seq_loop_monitor_4;
    seq_loop_intf#(276) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state17;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state21;
    assign seq_loop_intf_5.post_states_valid = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state20;
    assign seq_loop_intf_5.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_5.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state18;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state20;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(276) seq_loop_monitor_5;
    seq_loop_intf#(276) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state21;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state25;
    assign seq_loop_intf_6.post_states_valid = 1'b1;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state24;
    assign seq_loop_intf_6.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_6.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state22;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state24;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(276) seq_loop_monitor_6;
    seq_loop_intf#(276) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state25;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state29;
    assign seq_loop_intf_7.post_states_valid = 1'b1;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state28;
    assign seq_loop_intf_7.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_7.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state26;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state28;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(276) seq_loop_monitor_7;
    seq_loop_intf#(276) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state29;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state33;
    assign seq_loop_intf_8.post_states_valid = 1'b1;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state32;
    assign seq_loop_intf_8.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_8.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state30;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state32;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(276) seq_loop_monitor_8;
    seq_loop_intf#(276) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state33;
    assign seq_loop_intf_9.pre_states_valid = 1'b1;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state37;
    assign seq_loop_intf_9.post_states_valid = 1'b1;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state36;
    assign seq_loop_intf_9.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_9.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state34;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state36;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(276) seq_loop_monitor_9;
    seq_loop_intf#(276) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state37;
    assign seq_loop_intf_10.pre_states_valid = 1'b1;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state41;
    assign seq_loop_intf_10.post_states_valid = 1'b1;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state40;
    assign seq_loop_intf_10.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_10.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state38;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state40;
    assign seq_loop_intf_10.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(276) seq_loop_monitor_10;
    seq_loop_intf#(276) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state41;
    assign seq_loop_intf_11.pre_states_valid = 1'b1;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state45;
    assign seq_loop_intf_11.post_states_valid = 1'b1;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state44;
    assign seq_loop_intf_11.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_11.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state42;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state44;
    assign seq_loop_intf_11.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(276) seq_loop_monitor_11;
    seq_loop_intf#(276) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state45;
    assign seq_loop_intf_12.pre_states_valid = 1'b1;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state49;
    assign seq_loop_intf_12.post_states_valid = 1'b1;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state48;
    assign seq_loop_intf_12.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_12.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state46;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state48;
    assign seq_loop_intf_12.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(276) seq_loop_monitor_12;
    seq_loop_intf#(276) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state49;
    assign seq_loop_intf_13.pre_states_valid = 1'b1;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state53;
    assign seq_loop_intf_13.post_states_valid = 1'b1;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state52;
    assign seq_loop_intf_13.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_13.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state50;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state52;
    assign seq_loop_intf_13.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(276) seq_loop_monitor_13;
    seq_loop_intf#(276) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state53;
    assign seq_loop_intf_14.pre_states_valid = 1'b1;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state57;
    assign seq_loop_intf_14.post_states_valid = 1'b1;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state56;
    assign seq_loop_intf_14.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_14.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state54;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state56;
    assign seq_loop_intf_14.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(276) seq_loop_monitor_14;
    seq_loop_intf#(276) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state57;
    assign seq_loop_intf_15.pre_states_valid = 1'b1;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state61;
    assign seq_loop_intf_15.post_states_valid = 1'b1;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state60;
    assign seq_loop_intf_15.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_15.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state58;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state60;
    assign seq_loop_intf_15.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(276) seq_loop_monitor_15;
    seq_loop_intf#(276) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state61;
    assign seq_loop_intf_16.pre_states_valid = 1'b1;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state65;
    assign seq_loop_intf_16.post_states_valid = 1'b1;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state64;
    assign seq_loop_intf_16.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_16.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state62;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state64;
    assign seq_loop_intf_16.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(276) seq_loop_monitor_16;
    seq_loop_intf#(276) seq_loop_intf_17(clock,reset);
    assign seq_loop_intf_17.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state65;
    assign seq_loop_intf_17.pre_states_valid = 1'b1;
    assign seq_loop_intf_17.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state69;
    assign seq_loop_intf_17.post_states_valid = 1'b1;
    assign seq_loop_intf_17.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state68;
    assign seq_loop_intf_17.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_17.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_17.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state66;
    assign seq_loop_intf_17.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state68;
    assign seq_loop_intf_17.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_17.one_state_loop = 1'b0;
    assign seq_loop_intf_17.one_state_block = 1'b0;
    assign seq_loop_intf_17.finish = finish;
    csv_file_dump seq_loop_csv_dumper_17;
    seq_loop_monitor #(276) seq_loop_monitor_17;
    seq_loop_intf#(276) seq_loop_intf_18(clock,reset);
    assign seq_loop_intf_18.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state69;
    assign seq_loop_intf_18.pre_states_valid = 1'b1;
    assign seq_loop_intf_18.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state73;
    assign seq_loop_intf_18.post_states_valid = 1'b1;
    assign seq_loop_intf_18.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state72;
    assign seq_loop_intf_18.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_18.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_18.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state70;
    assign seq_loop_intf_18.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state72;
    assign seq_loop_intf_18.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_18.one_state_loop = 1'b0;
    assign seq_loop_intf_18.one_state_block = 1'b0;
    assign seq_loop_intf_18.finish = finish;
    csv_file_dump seq_loop_csv_dumper_18;
    seq_loop_monitor #(276) seq_loop_monitor_18;
    seq_loop_intf#(276) seq_loop_intf_19(clock,reset);
    assign seq_loop_intf_19.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state73;
    assign seq_loop_intf_19.pre_states_valid = 1'b1;
    assign seq_loop_intf_19.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state77;
    assign seq_loop_intf_19.post_states_valid = 1'b1;
    assign seq_loop_intf_19.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state76;
    assign seq_loop_intf_19.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_19.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_19.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state74;
    assign seq_loop_intf_19.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state76;
    assign seq_loop_intf_19.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_19.one_state_loop = 1'b0;
    assign seq_loop_intf_19.one_state_block = 1'b0;
    assign seq_loop_intf_19.finish = finish;
    csv_file_dump seq_loop_csv_dumper_19;
    seq_loop_monitor #(276) seq_loop_monitor_19;
    seq_loop_intf#(276) seq_loop_intf_20(clock,reset);
    assign seq_loop_intf_20.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state77;
    assign seq_loop_intf_20.pre_states_valid = 1'b1;
    assign seq_loop_intf_20.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state81;
    assign seq_loop_intf_20.post_states_valid = 1'b1;
    assign seq_loop_intf_20.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state80;
    assign seq_loop_intf_20.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_20.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_20.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state78;
    assign seq_loop_intf_20.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state80;
    assign seq_loop_intf_20.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_20.one_state_loop = 1'b0;
    assign seq_loop_intf_20.one_state_block = 1'b0;
    assign seq_loop_intf_20.finish = finish;
    csv_file_dump seq_loop_csv_dumper_20;
    seq_loop_monitor #(276) seq_loop_monitor_20;
    seq_loop_intf#(276) seq_loop_intf_21(clock,reset);
    assign seq_loop_intf_21.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state81;
    assign seq_loop_intf_21.pre_states_valid = 1'b1;
    assign seq_loop_intf_21.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state85;
    assign seq_loop_intf_21.post_states_valid = 1'b1;
    assign seq_loop_intf_21.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state84;
    assign seq_loop_intf_21.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_21.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_21.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state82;
    assign seq_loop_intf_21.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state84;
    assign seq_loop_intf_21.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_21.one_state_loop = 1'b0;
    assign seq_loop_intf_21.one_state_block = 1'b0;
    assign seq_loop_intf_21.finish = finish;
    csv_file_dump seq_loop_csv_dumper_21;
    seq_loop_monitor #(276) seq_loop_monitor_21;
    seq_loop_intf#(276) seq_loop_intf_22(clock,reset);
    assign seq_loop_intf_22.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state85;
    assign seq_loop_intf_22.pre_states_valid = 1'b1;
    assign seq_loop_intf_22.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state89;
    assign seq_loop_intf_22.post_states_valid = 1'b1;
    assign seq_loop_intf_22.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state88;
    assign seq_loop_intf_22.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_22.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_22.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_22.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state86;
    assign seq_loop_intf_22.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state88;
    assign seq_loop_intf_22.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_22.one_state_loop = 1'b0;
    assign seq_loop_intf_22.one_state_block = 1'b0;
    assign seq_loop_intf_22.finish = finish;
    csv_file_dump seq_loop_csv_dumper_22;
    seq_loop_monitor #(276) seq_loop_monitor_22;
    seq_loop_intf#(276) seq_loop_intf_23(clock,reset);
    assign seq_loop_intf_23.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state89;
    assign seq_loop_intf_23.pre_states_valid = 1'b1;
    assign seq_loop_intf_23.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state93;
    assign seq_loop_intf_23.post_states_valid = 1'b1;
    assign seq_loop_intf_23.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state92;
    assign seq_loop_intf_23.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_23.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_23.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state90;
    assign seq_loop_intf_23.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state92;
    assign seq_loop_intf_23.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_23.one_state_loop = 1'b0;
    assign seq_loop_intf_23.one_state_block = 1'b0;
    assign seq_loop_intf_23.finish = finish;
    csv_file_dump seq_loop_csv_dumper_23;
    seq_loop_monitor #(276) seq_loop_monitor_23;
    seq_loop_intf#(276) seq_loop_intf_24(clock,reset);
    assign seq_loop_intf_24.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state93;
    assign seq_loop_intf_24.pre_states_valid = 1'b1;
    assign seq_loop_intf_24.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state97;
    assign seq_loop_intf_24.post_states_valid = 1'b1;
    assign seq_loop_intf_24.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state96;
    assign seq_loop_intf_24.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_24.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_24.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state94;
    assign seq_loop_intf_24.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state96;
    assign seq_loop_intf_24.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_24.one_state_loop = 1'b0;
    assign seq_loop_intf_24.one_state_block = 1'b0;
    assign seq_loop_intf_24.finish = finish;
    csv_file_dump seq_loop_csv_dumper_24;
    seq_loop_monitor #(276) seq_loop_monitor_24;
    seq_loop_intf#(276) seq_loop_intf_25(clock,reset);
    assign seq_loop_intf_25.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state97;
    assign seq_loop_intf_25.pre_states_valid = 1'b1;
    assign seq_loop_intf_25.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state101;
    assign seq_loop_intf_25.post_states_valid = 1'b1;
    assign seq_loop_intf_25.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state100;
    assign seq_loop_intf_25.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_25.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_25.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state98;
    assign seq_loop_intf_25.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state100;
    assign seq_loop_intf_25.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_25.one_state_loop = 1'b0;
    assign seq_loop_intf_25.one_state_block = 1'b0;
    assign seq_loop_intf_25.finish = finish;
    csv_file_dump seq_loop_csv_dumper_25;
    seq_loop_monitor #(276) seq_loop_monitor_25;
    seq_loop_intf#(276) seq_loop_intf_26(clock,reset);
    assign seq_loop_intf_26.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state101;
    assign seq_loop_intf_26.pre_states_valid = 1'b1;
    assign seq_loop_intf_26.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state105;
    assign seq_loop_intf_26.post_states_valid = 1'b1;
    assign seq_loop_intf_26.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state104;
    assign seq_loop_intf_26.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_26.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_26.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state102;
    assign seq_loop_intf_26.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state104;
    assign seq_loop_intf_26.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_26.one_state_loop = 1'b0;
    assign seq_loop_intf_26.one_state_block = 1'b0;
    assign seq_loop_intf_26.finish = finish;
    csv_file_dump seq_loop_csv_dumper_26;
    seq_loop_monitor #(276) seq_loop_monitor_26;
    seq_loop_intf#(276) seq_loop_intf_27(clock,reset);
    assign seq_loop_intf_27.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state105;
    assign seq_loop_intf_27.pre_states_valid = 1'b1;
    assign seq_loop_intf_27.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state109;
    assign seq_loop_intf_27.post_states_valid = 1'b1;
    assign seq_loop_intf_27.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state108;
    assign seq_loop_intf_27.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_27.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_27.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state106;
    assign seq_loop_intf_27.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state108;
    assign seq_loop_intf_27.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_27.one_state_loop = 1'b0;
    assign seq_loop_intf_27.one_state_block = 1'b0;
    assign seq_loop_intf_27.finish = finish;
    csv_file_dump seq_loop_csv_dumper_27;
    seq_loop_monitor #(276) seq_loop_monitor_27;
    seq_loop_intf#(276) seq_loop_intf_28(clock,reset);
    assign seq_loop_intf_28.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state109;
    assign seq_loop_intf_28.pre_states_valid = 1'b1;
    assign seq_loop_intf_28.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state113;
    assign seq_loop_intf_28.post_states_valid = 1'b1;
    assign seq_loop_intf_28.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state112;
    assign seq_loop_intf_28.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_28.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_28.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state110;
    assign seq_loop_intf_28.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state112;
    assign seq_loop_intf_28.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_28.one_state_loop = 1'b0;
    assign seq_loop_intf_28.one_state_block = 1'b0;
    assign seq_loop_intf_28.finish = finish;
    csv_file_dump seq_loop_csv_dumper_28;
    seq_loop_monitor #(276) seq_loop_monitor_28;
    seq_loop_intf#(276) seq_loop_intf_29(clock,reset);
    assign seq_loop_intf_29.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state113;
    assign seq_loop_intf_29.pre_states_valid = 1'b1;
    assign seq_loop_intf_29.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state117;
    assign seq_loop_intf_29.post_states_valid = 1'b1;
    assign seq_loop_intf_29.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state116;
    assign seq_loop_intf_29.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_29.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_29.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state114;
    assign seq_loop_intf_29.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state116;
    assign seq_loop_intf_29.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_29.one_state_loop = 1'b0;
    assign seq_loop_intf_29.one_state_block = 1'b0;
    assign seq_loop_intf_29.finish = finish;
    csv_file_dump seq_loop_csv_dumper_29;
    seq_loop_monitor #(276) seq_loop_monitor_29;
    seq_loop_intf#(276) seq_loop_intf_30(clock,reset);
    assign seq_loop_intf_30.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state117;
    assign seq_loop_intf_30.pre_states_valid = 1'b1;
    assign seq_loop_intf_30.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state121;
    assign seq_loop_intf_30.post_states_valid = 1'b1;
    assign seq_loop_intf_30.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state120;
    assign seq_loop_intf_30.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_30.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_30.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state118;
    assign seq_loop_intf_30.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state120;
    assign seq_loop_intf_30.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_30.one_state_loop = 1'b0;
    assign seq_loop_intf_30.one_state_block = 1'b0;
    assign seq_loop_intf_30.finish = finish;
    csv_file_dump seq_loop_csv_dumper_30;
    seq_loop_monitor #(276) seq_loop_monitor_30;
    seq_loop_intf#(276) seq_loop_intf_31(clock,reset);
    assign seq_loop_intf_31.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state121;
    assign seq_loop_intf_31.pre_states_valid = 1'b1;
    assign seq_loop_intf_31.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state125;
    assign seq_loop_intf_31.post_states_valid = 1'b1;
    assign seq_loop_intf_31.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state124;
    assign seq_loop_intf_31.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_31.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_31.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state122;
    assign seq_loop_intf_31.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state124;
    assign seq_loop_intf_31.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_31.one_state_loop = 1'b0;
    assign seq_loop_intf_31.one_state_block = 1'b0;
    assign seq_loop_intf_31.finish = finish;
    csv_file_dump seq_loop_csv_dumper_31;
    seq_loop_monitor #(276) seq_loop_monitor_31;
    seq_loop_intf#(276) seq_loop_intf_32(clock,reset);
    assign seq_loop_intf_32.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state125;
    assign seq_loop_intf_32.pre_states_valid = 1'b1;
    assign seq_loop_intf_32.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state129;
    assign seq_loop_intf_32.post_states_valid = 1'b1;
    assign seq_loop_intf_32.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state128;
    assign seq_loop_intf_32.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_32.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_32.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state126;
    assign seq_loop_intf_32.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state128;
    assign seq_loop_intf_32.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_32.one_state_loop = 1'b0;
    assign seq_loop_intf_32.one_state_block = 1'b0;
    assign seq_loop_intf_32.finish = finish;
    csv_file_dump seq_loop_csv_dumper_32;
    seq_loop_monitor #(276) seq_loop_monitor_32;
    seq_loop_intf#(276) seq_loop_intf_33(clock,reset);
    assign seq_loop_intf_33.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state129;
    assign seq_loop_intf_33.pre_states_valid = 1'b1;
    assign seq_loop_intf_33.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state133;
    assign seq_loop_intf_33.post_states_valid = 1'b1;
    assign seq_loop_intf_33.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state132;
    assign seq_loop_intf_33.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_33.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_33.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state130;
    assign seq_loop_intf_33.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state132;
    assign seq_loop_intf_33.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_33.one_state_loop = 1'b0;
    assign seq_loop_intf_33.one_state_block = 1'b0;
    assign seq_loop_intf_33.finish = finish;
    csv_file_dump seq_loop_csv_dumper_33;
    seq_loop_monitor #(276) seq_loop_monitor_33;
    seq_loop_intf#(276) seq_loop_intf_34(clock,reset);
    assign seq_loop_intf_34.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state133;
    assign seq_loop_intf_34.pre_states_valid = 1'b1;
    assign seq_loop_intf_34.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state137;
    assign seq_loop_intf_34.post_states_valid = 1'b1;
    assign seq_loop_intf_34.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state136;
    assign seq_loop_intf_34.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_34.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_34.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state134;
    assign seq_loop_intf_34.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state136;
    assign seq_loop_intf_34.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_34.one_state_loop = 1'b0;
    assign seq_loop_intf_34.one_state_block = 1'b0;
    assign seq_loop_intf_34.finish = finish;
    csv_file_dump seq_loop_csv_dumper_34;
    seq_loop_monitor #(276) seq_loop_monitor_34;
    seq_loop_intf#(276) seq_loop_intf_35(clock,reset);
    assign seq_loop_intf_35.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state137;
    assign seq_loop_intf_35.pre_states_valid = 1'b1;
    assign seq_loop_intf_35.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state141;
    assign seq_loop_intf_35.post_states_valid = 1'b1;
    assign seq_loop_intf_35.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state140;
    assign seq_loop_intf_35.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_35.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_35.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state138;
    assign seq_loop_intf_35.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state140;
    assign seq_loop_intf_35.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_35.one_state_loop = 1'b0;
    assign seq_loop_intf_35.one_state_block = 1'b0;
    assign seq_loop_intf_35.finish = finish;
    csv_file_dump seq_loop_csv_dumper_35;
    seq_loop_monitor #(276) seq_loop_monitor_35;
    seq_loop_intf#(276) seq_loop_intf_36(clock,reset);
    assign seq_loop_intf_36.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state141;
    assign seq_loop_intf_36.pre_states_valid = 1'b1;
    assign seq_loop_intf_36.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state145;
    assign seq_loop_intf_36.post_states_valid = 1'b1;
    assign seq_loop_intf_36.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state144;
    assign seq_loop_intf_36.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_36.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_36.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_36.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_36.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state142;
    assign seq_loop_intf_36.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state144;
    assign seq_loop_intf_36.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_36.one_state_loop = 1'b0;
    assign seq_loop_intf_36.one_state_block = 1'b0;
    assign seq_loop_intf_36.finish = finish;
    csv_file_dump seq_loop_csv_dumper_36;
    seq_loop_monitor #(276) seq_loop_monitor_36;
    seq_loop_intf#(276) seq_loop_intf_37(clock,reset);
    assign seq_loop_intf_37.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state145;
    assign seq_loop_intf_37.pre_states_valid = 1'b1;
    assign seq_loop_intf_37.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state149;
    assign seq_loop_intf_37.post_states_valid = 1'b1;
    assign seq_loop_intf_37.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state148;
    assign seq_loop_intf_37.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_37.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_37.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_37.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_37.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state146;
    assign seq_loop_intf_37.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state148;
    assign seq_loop_intf_37.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_37.one_state_loop = 1'b0;
    assign seq_loop_intf_37.one_state_block = 1'b0;
    assign seq_loop_intf_37.finish = finish;
    csv_file_dump seq_loop_csv_dumper_37;
    seq_loop_monitor #(276) seq_loop_monitor_37;
    seq_loop_intf#(276) seq_loop_intf_38(clock,reset);
    assign seq_loop_intf_38.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state149;
    assign seq_loop_intf_38.pre_states_valid = 1'b1;
    assign seq_loop_intf_38.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state153;
    assign seq_loop_intf_38.post_states_valid = 1'b1;
    assign seq_loop_intf_38.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state152;
    assign seq_loop_intf_38.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_38.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_38.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_38.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_38.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state150;
    assign seq_loop_intf_38.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state152;
    assign seq_loop_intf_38.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_38.one_state_loop = 1'b0;
    assign seq_loop_intf_38.one_state_block = 1'b0;
    assign seq_loop_intf_38.finish = finish;
    csv_file_dump seq_loop_csv_dumper_38;
    seq_loop_monitor #(276) seq_loop_monitor_38;
    seq_loop_intf#(276) seq_loop_intf_39(clock,reset);
    assign seq_loop_intf_39.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state153;
    assign seq_loop_intf_39.pre_states_valid = 1'b1;
    assign seq_loop_intf_39.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state157;
    assign seq_loop_intf_39.post_states_valid = 1'b1;
    assign seq_loop_intf_39.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state156;
    assign seq_loop_intf_39.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_39.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_39.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_39.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_39.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state154;
    assign seq_loop_intf_39.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state156;
    assign seq_loop_intf_39.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_39.one_state_loop = 1'b0;
    assign seq_loop_intf_39.one_state_block = 1'b0;
    assign seq_loop_intf_39.finish = finish;
    csv_file_dump seq_loop_csv_dumper_39;
    seq_loop_monitor #(276) seq_loop_monitor_39;
    seq_loop_intf#(276) seq_loop_intf_40(clock,reset);
    assign seq_loop_intf_40.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state157;
    assign seq_loop_intf_40.pre_states_valid = 1'b1;
    assign seq_loop_intf_40.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state161;
    assign seq_loop_intf_40.post_states_valid = 1'b1;
    assign seq_loop_intf_40.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state160;
    assign seq_loop_intf_40.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_40.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_40.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_40.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_40.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state158;
    assign seq_loop_intf_40.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state160;
    assign seq_loop_intf_40.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_40.one_state_loop = 1'b0;
    assign seq_loop_intf_40.one_state_block = 1'b0;
    assign seq_loop_intf_40.finish = finish;
    csv_file_dump seq_loop_csv_dumper_40;
    seq_loop_monitor #(276) seq_loop_monitor_40;
    seq_loop_intf#(276) seq_loop_intf_41(clock,reset);
    assign seq_loop_intf_41.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state161;
    assign seq_loop_intf_41.pre_states_valid = 1'b1;
    assign seq_loop_intf_41.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state165;
    assign seq_loop_intf_41.post_states_valid = 1'b1;
    assign seq_loop_intf_41.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state164;
    assign seq_loop_intf_41.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_41.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_41.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_41.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_41.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state162;
    assign seq_loop_intf_41.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state164;
    assign seq_loop_intf_41.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_41.one_state_loop = 1'b0;
    assign seq_loop_intf_41.one_state_block = 1'b0;
    assign seq_loop_intf_41.finish = finish;
    csv_file_dump seq_loop_csv_dumper_41;
    seq_loop_monitor #(276) seq_loop_monitor_41;
    seq_loop_intf#(276) seq_loop_intf_42(clock,reset);
    assign seq_loop_intf_42.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state165;
    assign seq_loop_intf_42.pre_states_valid = 1'b1;
    assign seq_loop_intf_42.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state169;
    assign seq_loop_intf_42.post_states_valid = 1'b1;
    assign seq_loop_intf_42.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state168;
    assign seq_loop_intf_42.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_42.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_42.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_42.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_42.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state166;
    assign seq_loop_intf_42.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state168;
    assign seq_loop_intf_42.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_42.one_state_loop = 1'b0;
    assign seq_loop_intf_42.one_state_block = 1'b0;
    assign seq_loop_intf_42.finish = finish;
    csv_file_dump seq_loop_csv_dumper_42;
    seq_loop_monitor #(276) seq_loop_monitor_42;
    seq_loop_intf#(276) seq_loop_intf_43(clock,reset);
    assign seq_loop_intf_43.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state169;
    assign seq_loop_intf_43.pre_states_valid = 1'b1;
    assign seq_loop_intf_43.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state173;
    assign seq_loop_intf_43.post_states_valid = 1'b1;
    assign seq_loop_intf_43.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state172;
    assign seq_loop_intf_43.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_43.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_43.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_43.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_43.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state170;
    assign seq_loop_intf_43.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state172;
    assign seq_loop_intf_43.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_43.one_state_loop = 1'b0;
    assign seq_loop_intf_43.one_state_block = 1'b0;
    assign seq_loop_intf_43.finish = finish;
    csv_file_dump seq_loop_csv_dumper_43;
    seq_loop_monitor #(276) seq_loop_monitor_43;
    seq_loop_intf#(276) seq_loop_intf_44(clock,reset);
    assign seq_loop_intf_44.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state173;
    assign seq_loop_intf_44.pre_states_valid = 1'b1;
    assign seq_loop_intf_44.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state177;
    assign seq_loop_intf_44.post_states_valid = 1'b1;
    assign seq_loop_intf_44.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state176;
    assign seq_loop_intf_44.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_44.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_44.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_44.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_44.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state174;
    assign seq_loop_intf_44.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state176;
    assign seq_loop_intf_44.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_44.one_state_loop = 1'b0;
    assign seq_loop_intf_44.one_state_block = 1'b0;
    assign seq_loop_intf_44.finish = finish;
    csv_file_dump seq_loop_csv_dumper_44;
    seq_loop_monitor #(276) seq_loop_monitor_44;
    seq_loop_intf#(276) seq_loop_intf_45(clock,reset);
    assign seq_loop_intf_45.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state177;
    assign seq_loop_intf_45.pre_states_valid = 1'b1;
    assign seq_loop_intf_45.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state181;
    assign seq_loop_intf_45.post_states_valid = 1'b1;
    assign seq_loop_intf_45.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state180;
    assign seq_loop_intf_45.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_45.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_45.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_45.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_45.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state178;
    assign seq_loop_intf_45.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state180;
    assign seq_loop_intf_45.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_45.one_state_loop = 1'b0;
    assign seq_loop_intf_45.one_state_block = 1'b0;
    assign seq_loop_intf_45.finish = finish;
    csv_file_dump seq_loop_csv_dumper_45;
    seq_loop_monitor #(276) seq_loop_monitor_45;
    seq_loop_intf#(276) seq_loop_intf_46(clock,reset);
    assign seq_loop_intf_46.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state181;
    assign seq_loop_intf_46.pre_states_valid = 1'b1;
    assign seq_loop_intf_46.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state185;
    assign seq_loop_intf_46.post_states_valid = 1'b1;
    assign seq_loop_intf_46.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state184;
    assign seq_loop_intf_46.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_46.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_46.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_46.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_46.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state182;
    assign seq_loop_intf_46.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state184;
    assign seq_loop_intf_46.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_46.one_state_loop = 1'b0;
    assign seq_loop_intf_46.one_state_block = 1'b0;
    assign seq_loop_intf_46.finish = finish;
    csv_file_dump seq_loop_csv_dumper_46;
    seq_loop_monitor #(276) seq_loop_monitor_46;
    seq_loop_intf#(276) seq_loop_intf_47(clock,reset);
    assign seq_loop_intf_47.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state185;
    assign seq_loop_intf_47.pre_states_valid = 1'b1;
    assign seq_loop_intf_47.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state189;
    assign seq_loop_intf_47.post_states_valid = 1'b1;
    assign seq_loop_intf_47.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state188;
    assign seq_loop_intf_47.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_47.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_47.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_47.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_47.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state186;
    assign seq_loop_intf_47.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state188;
    assign seq_loop_intf_47.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_47.one_state_loop = 1'b0;
    assign seq_loop_intf_47.one_state_block = 1'b0;
    assign seq_loop_intf_47.finish = finish;
    csv_file_dump seq_loop_csv_dumper_47;
    seq_loop_monitor #(276) seq_loop_monitor_47;
    seq_loop_intf#(276) seq_loop_intf_48(clock,reset);
    assign seq_loop_intf_48.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state189;
    assign seq_loop_intf_48.pre_states_valid = 1'b1;
    assign seq_loop_intf_48.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state193;
    assign seq_loop_intf_48.post_states_valid = 1'b1;
    assign seq_loop_intf_48.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state192;
    assign seq_loop_intf_48.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_48.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_48.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_48.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_48.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state190;
    assign seq_loop_intf_48.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state192;
    assign seq_loop_intf_48.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_48.one_state_loop = 1'b0;
    assign seq_loop_intf_48.one_state_block = 1'b0;
    assign seq_loop_intf_48.finish = finish;
    csv_file_dump seq_loop_csv_dumper_48;
    seq_loop_monitor #(276) seq_loop_monitor_48;
    seq_loop_intf#(276) seq_loop_intf_49(clock,reset);
    assign seq_loop_intf_49.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state193;
    assign seq_loop_intf_49.pre_states_valid = 1'b1;
    assign seq_loop_intf_49.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state197;
    assign seq_loop_intf_49.post_states_valid = 1'b1;
    assign seq_loop_intf_49.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state196;
    assign seq_loop_intf_49.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_49.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_49.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_49.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_49.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state194;
    assign seq_loop_intf_49.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state196;
    assign seq_loop_intf_49.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_49.one_state_loop = 1'b0;
    assign seq_loop_intf_49.one_state_block = 1'b0;
    assign seq_loop_intf_49.finish = finish;
    csv_file_dump seq_loop_csv_dumper_49;
    seq_loop_monitor #(276) seq_loop_monitor_49;
    seq_loop_intf#(276) seq_loop_intf_50(clock,reset);
    assign seq_loop_intf_50.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state197;
    assign seq_loop_intf_50.pre_states_valid = 1'b1;
    assign seq_loop_intf_50.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state201;
    assign seq_loop_intf_50.post_states_valid = 1'b1;
    assign seq_loop_intf_50.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state200;
    assign seq_loop_intf_50.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_50.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_50.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_50.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_50.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state198;
    assign seq_loop_intf_50.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state200;
    assign seq_loop_intf_50.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_50.one_state_loop = 1'b0;
    assign seq_loop_intf_50.one_state_block = 1'b0;
    assign seq_loop_intf_50.finish = finish;
    csv_file_dump seq_loop_csv_dumper_50;
    seq_loop_monitor #(276) seq_loop_monitor_50;
    seq_loop_intf#(276) seq_loop_intf_51(clock,reset);
    assign seq_loop_intf_51.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state201;
    assign seq_loop_intf_51.pre_states_valid = 1'b1;
    assign seq_loop_intf_51.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state205;
    assign seq_loop_intf_51.post_states_valid = 1'b1;
    assign seq_loop_intf_51.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state204;
    assign seq_loop_intf_51.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_51.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_51.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_51.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_51.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state202;
    assign seq_loop_intf_51.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state204;
    assign seq_loop_intf_51.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_51.one_state_loop = 1'b0;
    assign seq_loop_intf_51.one_state_block = 1'b0;
    assign seq_loop_intf_51.finish = finish;
    csv_file_dump seq_loop_csv_dumper_51;
    seq_loop_monitor #(276) seq_loop_monitor_51;
    seq_loop_intf#(276) seq_loop_intf_52(clock,reset);
    assign seq_loop_intf_52.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state205;
    assign seq_loop_intf_52.pre_states_valid = 1'b1;
    assign seq_loop_intf_52.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state209;
    assign seq_loop_intf_52.post_states_valid = 1'b1;
    assign seq_loop_intf_52.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state208;
    assign seq_loop_intf_52.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_52.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_52.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_52.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_52.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state206;
    assign seq_loop_intf_52.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state208;
    assign seq_loop_intf_52.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_52.one_state_loop = 1'b0;
    assign seq_loop_intf_52.one_state_block = 1'b0;
    assign seq_loop_intf_52.finish = finish;
    csv_file_dump seq_loop_csv_dumper_52;
    seq_loop_monitor #(276) seq_loop_monitor_52;
    seq_loop_intf#(276) seq_loop_intf_53(clock,reset);
    assign seq_loop_intf_53.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state209;
    assign seq_loop_intf_53.pre_states_valid = 1'b1;
    assign seq_loop_intf_53.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state213;
    assign seq_loop_intf_53.post_states_valid = 1'b1;
    assign seq_loop_intf_53.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state212;
    assign seq_loop_intf_53.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_53.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_53.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_53.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_53.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state210;
    assign seq_loop_intf_53.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state212;
    assign seq_loop_intf_53.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_53.one_state_loop = 1'b0;
    assign seq_loop_intf_53.one_state_block = 1'b0;
    assign seq_loop_intf_53.finish = finish;
    csv_file_dump seq_loop_csv_dumper_53;
    seq_loop_monitor #(276) seq_loop_monitor_53;
    seq_loop_intf#(276) seq_loop_intf_54(clock,reset);
    assign seq_loop_intf_54.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state213;
    assign seq_loop_intf_54.pre_states_valid = 1'b1;
    assign seq_loop_intf_54.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state217;
    assign seq_loop_intf_54.post_states_valid = 1'b1;
    assign seq_loop_intf_54.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state216;
    assign seq_loop_intf_54.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_54.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_54.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_54.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_54.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state214;
    assign seq_loop_intf_54.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state216;
    assign seq_loop_intf_54.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_54.one_state_loop = 1'b0;
    assign seq_loop_intf_54.one_state_block = 1'b0;
    assign seq_loop_intf_54.finish = finish;
    csv_file_dump seq_loop_csv_dumper_54;
    seq_loop_monitor #(276) seq_loop_monitor_54;
    seq_loop_intf#(276) seq_loop_intf_55(clock,reset);
    assign seq_loop_intf_55.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state217;
    assign seq_loop_intf_55.pre_states_valid = 1'b1;
    assign seq_loop_intf_55.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state221;
    assign seq_loop_intf_55.post_states_valid = 1'b1;
    assign seq_loop_intf_55.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state220;
    assign seq_loop_intf_55.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_55.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_55.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_55.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_55.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state218;
    assign seq_loop_intf_55.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state220;
    assign seq_loop_intf_55.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_55.one_state_loop = 1'b0;
    assign seq_loop_intf_55.one_state_block = 1'b0;
    assign seq_loop_intf_55.finish = finish;
    csv_file_dump seq_loop_csv_dumper_55;
    seq_loop_monitor #(276) seq_loop_monitor_55;
    seq_loop_intf#(276) seq_loop_intf_56(clock,reset);
    assign seq_loop_intf_56.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state221;
    assign seq_loop_intf_56.pre_states_valid = 1'b1;
    assign seq_loop_intf_56.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state225;
    assign seq_loop_intf_56.post_states_valid = 1'b1;
    assign seq_loop_intf_56.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state224;
    assign seq_loop_intf_56.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_56.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_56.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_56.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_56.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state222;
    assign seq_loop_intf_56.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state224;
    assign seq_loop_intf_56.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_56.one_state_loop = 1'b0;
    assign seq_loop_intf_56.one_state_block = 1'b0;
    assign seq_loop_intf_56.finish = finish;
    csv_file_dump seq_loop_csv_dumper_56;
    seq_loop_monitor #(276) seq_loop_monitor_56;
    seq_loop_intf#(276) seq_loop_intf_57(clock,reset);
    assign seq_loop_intf_57.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state225;
    assign seq_loop_intf_57.pre_states_valid = 1'b1;
    assign seq_loop_intf_57.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state229;
    assign seq_loop_intf_57.post_states_valid = 1'b1;
    assign seq_loop_intf_57.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state228;
    assign seq_loop_intf_57.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_57.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_57.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_57.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_57.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state226;
    assign seq_loop_intf_57.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state228;
    assign seq_loop_intf_57.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_57.one_state_loop = 1'b0;
    assign seq_loop_intf_57.one_state_block = 1'b0;
    assign seq_loop_intf_57.finish = finish;
    csv_file_dump seq_loop_csv_dumper_57;
    seq_loop_monitor #(276) seq_loop_monitor_57;
    seq_loop_intf#(276) seq_loop_intf_58(clock,reset);
    assign seq_loop_intf_58.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state229;
    assign seq_loop_intf_58.pre_states_valid = 1'b1;
    assign seq_loop_intf_58.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state233;
    assign seq_loop_intf_58.post_states_valid = 1'b1;
    assign seq_loop_intf_58.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state232;
    assign seq_loop_intf_58.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_58.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_58.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_58.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_58.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state230;
    assign seq_loop_intf_58.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state232;
    assign seq_loop_intf_58.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_58.one_state_loop = 1'b0;
    assign seq_loop_intf_58.one_state_block = 1'b0;
    assign seq_loop_intf_58.finish = finish;
    csv_file_dump seq_loop_csv_dumper_58;
    seq_loop_monitor #(276) seq_loop_monitor_58;
    seq_loop_intf#(276) seq_loop_intf_59(clock,reset);
    assign seq_loop_intf_59.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state233;
    assign seq_loop_intf_59.pre_states_valid = 1'b1;
    assign seq_loop_intf_59.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state237;
    assign seq_loop_intf_59.post_states_valid = 1'b1;
    assign seq_loop_intf_59.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state236;
    assign seq_loop_intf_59.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_59.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_59.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_59.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_59.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state234;
    assign seq_loop_intf_59.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state236;
    assign seq_loop_intf_59.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_59.one_state_loop = 1'b0;
    assign seq_loop_intf_59.one_state_block = 1'b0;
    assign seq_loop_intf_59.finish = finish;
    csv_file_dump seq_loop_csv_dumper_59;
    seq_loop_monitor #(276) seq_loop_monitor_59;
    seq_loop_intf#(276) seq_loop_intf_60(clock,reset);
    assign seq_loop_intf_60.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state237;
    assign seq_loop_intf_60.pre_states_valid = 1'b1;
    assign seq_loop_intf_60.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state241;
    assign seq_loop_intf_60.post_states_valid = 1'b1;
    assign seq_loop_intf_60.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state240;
    assign seq_loop_intf_60.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_60.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_60.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_60.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_60.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state238;
    assign seq_loop_intf_60.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state240;
    assign seq_loop_intf_60.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_60.one_state_loop = 1'b0;
    assign seq_loop_intf_60.one_state_block = 1'b0;
    assign seq_loop_intf_60.finish = finish;
    csv_file_dump seq_loop_csv_dumper_60;
    seq_loop_monitor #(276) seq_loop_monitor_60;
    seq_loop_intf#(276) seq_loop_intf_61(clock,reset);
    assign seq_loop_intf_61.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state241;
    assign seq_loop_intf_61.pre_states_valid = 1'b1;
    assign seq_loop_intf_61.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state245;
    assign seq_loop_intf_61.post_states_valid = 1'b1;
    assign seq_loop_intf_61.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state244;
    assign seq_loop_intf_61.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_61.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_61.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_61.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_61.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state242;
    assign seq_loop_intf_61.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state244;
    assign seq_loop_intf_61.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_61.one_state_loop = 1'b0;
    assign seq_loop_intf_61.one_state_block = 1'b0;
    assign seq_loop_intf_61.finish = finish;
    csv_file_dump seq_loop_csv_dumper_61;
    seq_loop_monitor #(276) seq_loop_monitor_61;
    seq_loop_intf#(276) seq_loop_intf_62(clock,reset);
    assign seq_loop_intf_62.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state245;
    assign seq_loop_intf_62.pre_states_valid = 1'b1;
    assign seq_loop_intf_62.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state249;
    assign seq_loop_intf_62.post_states_valid = 1'b1;
    assign seq_loop_intf_62.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state248;
    assign seq_loop_intf_62.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_62.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_62.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_62.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_62.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state246;
    assign seq_loop_intf_62.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state248;
    assign seq_loop_intf_62.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_62.one_state_loop = 1'b0;
    assign seq_loop_intf_62.one_state_block = 1'b0;
    assign seq_loop_intf_62.finish = finish;
    csv_file_dump seq_loop_csv_dumper_62;
    seq_loop_monitor #(276) seq_loop_monitor_62;
    seq_loop_intf#(276) seq_loop_intf_63(clock,reset);
    assign seq_loop_intf_63.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state249;
    assign seq_loop_intf_63.pre_states_valid = 1'b1;
    assign seq_loop_intf_63.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state253;
    assign seq_loop_intf_63.post_states_valid = 1'b1;
    assign seq_loop_intf_63.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state252;
    assign seq_loop_intf_63.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_63.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_63.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_63.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_63.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state250;
    assign seq_loop_intf_63.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state252;
    assign seq_loop_intf_63.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_63.one_state_loop = 1'b0;
    assign seq_loop_intf_63.one_state_block = 1'b0;
    assign seq_loop_intf_63.finish = finish;
    csv_file_dump seq_loop_csv_dumper_63;
    seq_loop_monitor #(276) seq_loop_monitor_63;
    seq_loop_intf#(276) seq_loop_intf_64(clock,reset);
    assign seq_loop_intf_64.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state253;
    assign seq_loop_intf_64.pre_states_valid = 1'b1;
    assign seq_loop_intf_64.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state257;
    assign seq_loop_intf_64.post_states_valid = 1'b1;
    assign seq_loop_intf_64.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state256;
    assign seq_loop_intf_64.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_64.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_64.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_64.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_64.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state254;
    assign seq_loop_intf_64.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state256;
    assign seq_loop_intf_64.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_64.one_state_loop = 1'b0;
    assign seq_loop_intf_64.one_state_block = 1'b0;
    assign seq_loop_intf_64.finish = finish;
    csv_file_dump seq_loop_csv_dumper_64;
    seq_loop_monitor #(276) seq_loop_monitor_64;
    seq_loop_intf#(276) seq_loop_intf_65(clock,reset);
    assign seq_loop_intf_65.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state257;
    assign seq_loop_intf_65.pre_states_valid = 1'b1;
    assign seq_loop_intf_65.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state261;
    assign seq_loop_intf_65.post_states_valid = 1'b1;
    assign seq_loop_intf_65.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state260;
    assign seq_loop_intf_65.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_65.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_65.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_65.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_65.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state258;
    assign seq_loop_intf_65.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state260;
    assign seq_loop_intf_65.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_65.one_state_loop = 1'b0;
    assign seq_loop_intf_65.one_state_block = 1'b0;
    assign seq_loop_intf_65.finish = finish;
    csv_file_dump seq_loop_csv_dumper_65;
    seq_loop_monitor #(276) seq_loop_monitor_65;
    seq_loop_intf#(276) seq_loop_intf_66(clock,reset);
    assign seq_loop_intf_66.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state3;
    assign seq_loop_intf_66.pre_states_valid = 1'b1;
    assign seq_loop_intf_66.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state270;
    assign seq_loop_intf_66.post_states_valid = 1'b1;
    assign seq_loop_intf_66.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state4;
    assign seq_loop_intf_66.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_66.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_66.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_66.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_66.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state4;
    assign seq_loop_intf_66.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state261;
    assign seq_loop_intf_66.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_66.one_state_loop = 1'b0;
    assign seq_loop_intf_66.one_state_block = 1'b0;
    assign seq_loop_intf_66.finish = finish;
    csv_file_dump seq_loop_csv_dumper_66;
    seq_loop_monitor #(276) seq_loop_monitor_66;
    seq_loop_intf#(276) seq_loop_intf_67(clock,reset);
    assign seq_loop_intf_67.pre_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state270;
    assign seq_loop_intf_67.pre_states_valid = 1'b1;
    assign seq_loop_intf_67.post_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state276;
    assign seq_loop_intf_67.post_states_valid = 1'b1;
    assign seq_loop_intf_67.quit_loop_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state271;
    assign seq_loop_intf_67.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_67.quit_loop_state1 = 276'h0;
    assign seq_loop_intf_67.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_67.cur_state = AESL_inst_test_state_buffer.ap_CS_fsm;
    assign seq_loop_intf_67.iter_start_state = AESL_inst_test_state_buffer.ap_ST_fsm_state271;
    assign seq_loop_intf_67.iter_end_state0 = AESL_inst_test_state_buffer.ap_ST_fsm_state275;
    assign seq_loop_intf_67.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_67.one_state_loop = 1'b0;
    assign seq_loop_intf_67.one_state_block = 1'b0;
    assign seq_loop_intf_67.finish = finish;
    csv_file_dump seq_loop_csv_dumper_67;
    seq_loop_monitor #(276) seq_loop_monitor_67;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.loop_start = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_test_state_buffer.grp_test_state_buffer_Pipeline_VITIS_LOOP_43_3_fu_7502.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b0;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);
    seq_loop_csv_dumper_17 = new("./seq_loop_status17.csv");
    seq_loop_monitor_17 = new(seq_loop_intf_17,seq_loop_csv_dumper_17);
    seq_loop_csv_dumper_18 = new("./seq_loop_status18.csv");
    seq_loop_monitor_18 = new(seq_loop_intf_18,seq_loop_csv_dumper_18);
    seq_loop_csv_dumper_19 = new("./seq_loop_status19.csv");
    seq_loop_monitor_19 = new(seq_loop_intf_19,seq_loop_csv_dumper_19);
    seq_loop_csv_dumper_20 = new("./seq_loop_status20.csv");
    seq_loop_monitor_20 = new(seq_loop_intf_20,seq_loop_csv_dumper_20);
    seq_loop_csv_dumper_21 = new("./seq_loop_status21.csv");
    seq_loop_monitor_21 = new(seq_loop_intf_21,seq_loop_csv_dumper_21);
    seq_loop_csv_dumper_22 = new("./seq_loop_status22.csv");
    seq_loop_monitor_22 = new(seq_loop_intf_22,seq_loop_csv_dumper_22);
    seq_loop_csv_dumper_23 = new("./seq_loop_status23.csv");
    seq_loop_monitor_23 = new(seq_loop_intf_23,seq_loop_csv_dumper_23);
    seq_loop_csv_dumper_24 = new("./seq_loop_status24.csv");
    seq_loop_monitor_24 = new(seq_loop_intf_24,seq_loop_csv_dumper_24);
    seq_loop_csv_dumper_25 = new("./seq_loop_status25.csv");
    seq_loop_monitor_25 = new(seq_loop_intf_25,seq_loop_csv_dumper_25);
    seq_loop_csv_dumper_26 = new("./seq_loop_status26.csv");
    seq_loop_monitor_26 = new(seq_loop_intf_26,seq_loop_csv_dumper_26);
    seq_loop_csv_dumper_27 = new("./seq_loop_status27.csv");
    seq_loop_monitor_27 = new(seq_loop_intf_27,seq_loop_csv_dumper_27);
    seq_loop_csv_dumper_28 = new("./seq_loop_status28.csv");
    seq_loop_monitor_28 = new(seq_loop_intf_28,seq_loop_csv_dumper_28);
    seq_loop_csv_dumper_29 = new("./seq_loop_status29.csv");
    seq_loop_monitor_29 = new(seq_loop_intf_29,seq_loop_csv_dumper_29);
    seq_loop_csv_dumper_30 = new("./seq_loop_status30.csv");
    seq_loop_monitor_30 = new(seq_loop_intf_30,seq_loop_csv_dumper_30);
    seq_loop_csv_dumper_31 = new("./seq_loop_status31.csv");
    seq_loop_monitor_31 = new(seq_loop_intf_31,seq_loop_csv_dumper_31);
    seq_loop_csv_dumper_32 = new("./seq_loop_status32.csv");
    seq_loop_monitor_32 = new(seq_loop_intf_32,seq_loop_csv_dumper_32);
    seq_loop_csv_dumper_33 = new("./seq_loop_status33.csv");
    seq_loop_monitor_33 = new(seq_loop_intf_33,seq_loop_csv_dumper_33);
    seq_loop_csv_dumper_34 = new("./seq_loop_status34.csv");
    seq_loop_monitor_34 = new(seq_loop_intf_34,seq_loop_csv_dumper_34);
    seq_loop_csv_dumper_35 = new("./seq_loop_status35.csv");
    seq_loop_monitor_35 = new(seq_loop_intf_35,seq_loop_csv_dumper_35);
    seq_loop_csv_dumper_36 = new("./seq_loop_status36.csv");
    seq_loop_monitor_36 = new(seq_loop_intf_36,seq_loop_csv_dumper_36);
    seq_loop_csv_dumper_37 = new("./seq_loop_status37.csv");
    seq_loop_monitor_37 = new(seq_loop_intf_37,seq_loop_csv_dumper_37);
    seq_loop_csv_dumper_38 = new("./seq_loop_status38.csv");
    seq_loop_monitor_38 = new(seq_loop_intf_38,seq_loop_csv_dumper_38);
    seq_loop_csv_dumper_39 = new("./seq_loop_status39.csv");
    seq_loop_monitor_39 = new(seq_loop_intf_39,seq_loop_csv_dumper_39);
    seq_loop_csv_dumper_40 = new("./seq_loop_status40.csv");
    seq_loop_monitor_40 = new(seq_loop_intf_40,seq_loop_csv_dumper_40);
    seq_loop_csv_dumper_41 = new("./seq_loop_status41.csv");
    seq_loop_monitor_41 = new(seq_loop_intf_41,seq_loop_csv_dumper_41);
    seq_loop_csv_dumper_42 = new("./seq_loop_status42.csv");
    seq_loop_monitor_42 = new(seq_loop_intf_42,seq_loop_csv_dumper_42);
    seq_loop_csv_dumper_43 = new("./seq_loop_status43.csv");
    seq_loop_monitor_43 = new(seq_loop_intf_43,seq_loop_csv_dumper_43);
    seq_loop_csv_dumper_44 = new("./seq_loop_status44.csv");
    seq_loop_monitor_44 = new(seq_loop_intf_44,seq_loop_csv_dumper_44);
    seq_loop_csv_dumper_45 = new("./seq_loop_status45.csv");
    seq_loop_monitor_45 = new(seq_loop_intf_45,seq_loop_csv_dumper_45);
    seq_loop_csv_dumper_46 = new("./seq_loop_status46.csv");
    seq_loop_monitor_46 = new(seq_loop_intf_46,seq_loop_csv_dumper_46);
    seq_loop_csv_dumper_47 = new("./seq_loop_status47.csv");
    seq_loop_monitor_47 = new(seq_loop_intf_47,seq_loop_csv_dumper_47);
    seq_loop_csv_dumper_48 = new("./seq_loop_status48.csv");
    seq_loop_monitor_48 = new(seq_loop_intf_48,seq_loop_csv_dumper_48);
    seq_loop_csv_dumper_49 = new("./seq_loop_status49.csv");
    seq_loop_monitor_49 = new(seq_loop_intf_49,seq_loop_csv_dumper_49);
    seq_loop_csv_dumper_50 = new("./seq_loop_status50.csv");
    seq_loop_monitor_50 = new(seq_loop_intf_50,seq_loop_csv_dumper_50);
    seq_loop_csv_dumper_51 = new("./seq_loop_status51.csv");
    seq_loop_monitor_51 = new(seq_loop_intf_51,seq_loop_csv_dumper_51);
    seq_loop_csv_dumper_52 = new("./seq_loop_status52.csv");
    seq_loop_monitor_52 = new(seq_loop_intf_52,seq_loop_csv_dumper_52);
    seq_loop_csv_dumper_53 = new("./seq_loop_status53.csv");
    seq_loop_monitor_53 = new(seq_loop_intf_53,seq_loop_csv_dumper_53);
    seq_loop_csv_dumper_54 = new("./seq_loop_status54.csv");
    seq_loop_monitor_54 = new(seq_loop_intf_54,seq_loop_csv_dumper_54);
    seq_loop_csv_dumper_55 = new("./seq_loop_status55.csv");
    seq_loop_monitor_55 = new(seq_loop_intf_55,seq_loop_csv_dumper_55);
    seq_loop_csv_dumper_56 = new("./seq_loop_status56.csv");
    seq_loop_monitor_56 = new(seq_loop_intf_56,seq_loop_csv_dumper_56);
    seq_loop_csv_dumper_57 = new("./seq_loop_status57.csv");
    seq_loop_monitor_57 = new(seq_loop_intf_57,seq_loop_csv_dumper_57);
    seq_loop_csv_dumper_58 = new("./seq_loop_status58.csv");
    seq_loop_monitor_58 = new(seq_loop_intf_58,seq_loop_csv_dumper_58);
    seq_loop_csv_dumper_59 = new("./seq_loop_status59.csv");
    seq_loop_monitor_59 = new(seq_loop_intf_59,seq_loop_csv_dumper_59);
    seq_loop_csv_dumper_60 = new("./seq_loop_status60.csv");
    seq_loop_monitor_60 = new(seq_loop_intf_60,seq_loop_csv_dumper_60);
    seq_loop_csv_dumper_61 = new("./seq_loop_status61.csv");
    seq_loop_monitor_61 = new(seq_loop_intf_61,seq_loop_csv_dumper_61);
    seq_loop_csv_dumper_62 = new("./seq_loop_status62.csv");
    seq_loop_monitor_62 = new(seq_loop_intf_62,seq_loop_csv_dumper_62);
    seq_loop_csv_dumper_63 = new("./seq_loop_status63.csv");
    seq_loop_monitor_63 = new(seq_loop_intf_63,seq_loop_csv_dumper_63);
    seq_loop_csv_dumper_64 = new("./seq_loop_status64.csv");
    seq_loop_monitor_64 = new(seq_loop_intf_64,seq_loop_csv_dumper_64);
    seq_loop_csv_dumper_65 = new("./seq_loop_status65.csv");
    seq_loop_monitor_65 = new(seq_loop_intf_65,seq_loop_csv_dumper_65);
    seq_loop_csv_dumper_66 = new("./seq_loop_status66.csv");
    seq_loop_monitor_66 = new(seq_loop_intf_66,seq_loop_csv_dumper_66);
    seq_loop_csv_dumper_67 = new("./seq_loop_status67.csv");
    seq_loop_monitor_67 = new(seq_loop_intf_67,seq_loop_csv_dumper_67);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_19);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_20);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_21);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_22);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_23);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_24);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_25);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_26);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_27);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_28);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_29);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_30);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_31);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_32);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_33);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_34);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_35);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_36);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_37);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_38);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_39);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_40);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_41);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_42);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_43);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_44);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_45);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_46);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_47);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_48);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_49);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_50);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_51);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_52);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_53);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_54);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_55);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_56);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_57);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_58);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_59);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_60);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_61);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_62);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_63);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_64);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_65);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_66);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_67);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
